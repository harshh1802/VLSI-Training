library verilog;
use verilog.vl_types.all;
entity ram_defines_sv_unit is
end ram_defines_sv_unit;
