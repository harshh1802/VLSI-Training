library verilog;
use verilog.vl_types.all;
entity ram_generator_sv_unit is
end ram_generator_sv_unit;
