library verilog;
use verilog.vl_types.all;
entity trans is
end trans;
