library verilog;
use verilog.vl_types.all;
entity ram_driver_sv_unit is
end ram_driver_sv_unit;
