library verilog;
use verilog.vl_types.all;
entity ram_trans_sv_unit is
end ram_trans_sv_unit;
