library verilog;
use verilog.vl_types.all;
entity ram_interface is
    port(
        clk             : in     vl_logic
    );
end ram_interface;
