class ram_base_test;

  //take handle of verification environment class
  
  //declare all interface 
  
   //take connect method (only for virtual interface)
   
   //create environment and call its methods here as needed
   function void build();
    :
   endtask
   
   function void connect(...);
    :
   endtask
   
   task run();
    :
   endtask
     
  
endclass